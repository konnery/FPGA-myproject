library verilog;
use verilog.vl_types.all;
entity da_tb is
end da_tb;
